
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY iir_IP IS
  PORT( clk                               :   IN    std_logic;
        reset                             :   IN    std_logic;
        clk_enable                        :   IN    std_logic;
        dataIn                            :   IN    std_logic_vector(15 DOWNTO 0);  -- sfix16_En8
        validIn                           :   IN    std_logic;
        ce_out                            :   OUT   std_logic;
        dataOut                           :   OUT   std_logic_vector(15 DOWNTO 0);  -- sfix16_En15
        validOut                          :   OUT   std_logic
        );
END iir_IP;


ARCHITECTURE rtl OF iir_IP IS

  -- Component Declarations
  COMPONENT dsphdl_BiquadFilter
    PORT( clk                             :   IN    std_logic;
          reset                           :   IN    std_logic;
          enb                             :   IN    std_logic;
          dataIn                          :   IN    std_logic_vector(15 DOWNTO 0);  -- sfix16_En8
          validIn                         :   IN    std_logic;
          dataOut                         :   OUT   std_logic_vector(15 DOWNTO 0);  -- sfix16_En15
          validOut                        :   OUT   std_logic
          );
  END COMPONENT;

  -- Component Configuration Statements
  FOR ALL : dsphdl_BiquadFilter
    USE ENTITY work.dsphdl_BiquadFilter(rtl);

  -- Signals
  SIGNAL varargout_1                      : std_logic_vector(15 DOWNTO 0);  -- ufix16
  SIGNAL varargout_2                      : std_logic;

BEGIN
  -- Generated by HDL IP Designer.
  u_dsphdl_BiquadFilter : dsphdl_BiquadFilter
    PORT MAP( clk => clk,
              reset => reset,
              enb => clk_enable,
              dataIn => dataIn,  -- sfix16_En8
              validIn => validIn,
              dataOut => varargout_1,  -- sfix16_En15
              validOut => varargout_2
              );

  ce_out <= clk_enable;

  dataOut <= varargout_1;

  validOut <= varargout_2;

END rtl;

